
module multiplier #(
    parameter N_IN = 4,
    parameter N_OUT = 8
    ) (
    input logic [N_IN-1:0] operand_a_i,
    input logic [N_IN-1:0] operand_b_i,
    output logic [N_OUT-1:0] result_o
);

assign result_o

endmodule
